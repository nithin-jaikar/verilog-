module basic(a,b,c);
	input a,c;
	output b;
	assign b = a && c ;
endmodule
	
